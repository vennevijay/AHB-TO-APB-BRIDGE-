class env_config extends uvm_object;
	`uvm_object_utils(env_config)

	int has_master_agent=1;
	int has_slave_agent=1;

	int no_of_master_agents=1;
	int no_of_slave_agents=1;

	int has_scoreboard=1;
	
	master_config m_cfg;
	slave_config s_cfg;

	extern function new(string name="env_config");	
		

endclass

	function env_config::new(string name);
		super.new(name);
	endfunction


